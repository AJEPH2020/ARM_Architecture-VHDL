library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;

entity dataMemory is
port(
    clk: in std_logic;
    writeOnDm: in std_logic;
    adrsdm: in std_logic_vector(5 downto 0);
    Din: in std_logic_vector(31 downto 0);
    bytes: in std_logic_vector(3 downto 0);
    outputdm: out std_logic_vector(31 downto 0);

    adrspm: IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    outputpm: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
    );
end entity;


architecture bev of dataMemory is

type mem is array(0 to 127) of std_logic_vector(31 downto 0);
signal add: integer range 0 to 127;

SIGNAL dmemory: mem:=(
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    
    X"E3A0100A",
    X"E3A02011",
    X"E0810002",
    X"E4810004",
    X"E1C100B0",
    X"E5E10005",
    X"E5913000",
    X"E1D140B0",
    X"E1D150F0",
    X"E5D16000",
    X"E1D170D0",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000",
    "00000000000000000000000000000000"
);


begin
	process(clk)
    begin
    	add<=conv_integer(adrsdm);
        outputdm<=dmemory(add);
        if(rising_edge(clk)) then
            if (writeOnDm = '1') then
                case bytes is
                    when "0001"=>
                        dmemory(add)(7 downto 0)<=Din(7 downto 0);
                    when "0010"=>
                        dmemory(add)(15 downto 8)<=Din(15 downto 8);
                    when "0011"=>
                        dmemory(add)(15 downto 0)<=Din(15 downto 0);
                    when "0100"=>
                        dmemory(add)(23 downto 16)<=Din(23 downto 16);
                    when "0101"=>
                        dmemory(add)(23 downto 16)<=Din(23 downto 16);
                        dmemory(add)(7 downto 0)<=Din(7 downto 0);
                    when "0110"=>
                        dmemory(add)(23 downto 8)<=Din(23 downto 8);
                    when "0111"=>
                        dmemory(add)(23 downto 0)<=Din(23 downto 0);
                    when "1000"=>
                        dmemory(add)(31 downto 24)<=Din(31 downto 24);
                    when "1001"=>
                        dmemory(add)(31 downto 24)<=Din(31 downto 24);
                        dmemory(add)(7 downto 0)<=Din(7 downto 0);
                    when "1010"=>
                        dmemory(add)(31 downto 24)<=Din(31 downto 24);
                        dmemory(add)(15 downto 8)<=Din(15 downto 8);
                    when "1011"=>
                        dmemory(add)(31 downto 24)<=Din(31 downto 24);
                        dmemory(add)(15 downto 0)<=Din(15 downto 0);
                    when "1100"=>
                        dmemory(add)(31 downto 16)<=Din(31 downto 16);
                    when "1101"=>
                        dmemory(add)(31 downto 16)<=Din(31 downto 16);
                        dmemory(add)(7 downto 0)<=Din(7 downto 0);
                    when "1110"=>
                        dmemory(add)(31 downto 8)<=Din(31 downto 8);
                    when "1111"=>
                        dmemory(add)<=Din;
                    when others=>
                        dmemory(add)<="ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";
                end case;
            end if;
        end if;

	end process;

    process(adrspm)
    begin
        outputpm<=dmemory(CONV_INTEGER(adrspm) + 64);
    end process;

end bev;

